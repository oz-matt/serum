package axil_if_c;
	`include "protocol_checker/axi_raddr_props.sv"
	`include "protocol_checker/axi_rdata_props.sv" 
	`include "protocol_checker/axi_waddr_props.sv"
	`include "protocol_checker/axi_wdata_props.sv"
	`include "protocol_checker/axi_wresp_props.sv"
endpackage